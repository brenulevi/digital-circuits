clock_counter_inst : clock_counter PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
