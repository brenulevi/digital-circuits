library ieee;
use ieee.std_logic_1164.all;

entity letter is
	port (
		KEY: 	in std_logic_vector(3 downto 0);
		SW: 	in std_logic_vector(9 downto 0);
		CLOCK_50 : in std_logic;
		HEX0: out std_logic_vector(6 downto 0);
		HEX1: out std_logic_vector(6 downto 0);
		HEX2: out std_logic_vector(6 downto 0);
		HEX3: out std_logic_vector(6 downto 0);
		LEDR:	out std_logic_vector(9 downto 0);
		LEDG: out std_logic_vector(7 downto 0)
	);
end entity letter;

architecture letter_arc of letter is

	component clock_counter is
		port (
			CLOCK_50 : in std_logic;
			CLOCK_4HZ : out std_logic
		);
	end component clock_counter;

	component mux is
		port (
			A,B, SEL: in std_logic;
			OTPT: out std_logic
		);
	end component mux;
	
	component counter is
		port (
			CLK, RST : in std_logic;
			OTPT : out std_logic_vector(3 downto 0)
		);
	end component counter;
	
	component adder is
		port (
			N : in std_logic_vector(3 downto 0);
			S : in std_logic_vector(3 downto 0);
			OTPT: out std_logic_vector(3 downto 0)
		);
	end component adder;
	
	component decodifier is
		port (
			A: in std_logic_vector(3 downto 0);
			OTPT: out std_logic_vector(6 downto 0)
		);
	end component decodifier;

	signal MUX_OTPT : std_logic;
	signal COUNTER_OTPT : std_logic_vector(3 downto 0);
	signal ADDER1_OTPT : std_logic_vector(3 downto 0);
	signal ADDER2_OTPT : std_logic_vector(3 downto 0);
	signal ADDER3_OTPT : std_logic_vector(3 downto 0);
	signal CLOCK_4HZ : std_logic;
	signal clk : std_logic;
begin

	-- 1 clock counter (made by Quartus Super Function) (Gets counter[23] to reduce the clock frequency) (actual = 4hz (i think))
	clock_counter1 : clock_counter port map (CLOCK_50 => CLOCK_50, CLOCK_4HZ => CLOCK_4HZ);
	
	-- 1 mux (selector between auto clock and manual clock based on switch (SW(0)))
	mux1: mux port map (A => not KEY(0), B => CLOCK_4HZ, SEL => SW(0), OTPT => MUX_OTPT);
	
	-- 1 instance of counter (0 to 7 | 4 bits)
	counter1 : counter port map (CLK => MUX_OTPT, RST => not KEY(3), OTPT => COUNTER_OTPT);

	-- 3 adder (counter + 1, counter + 2, counter + 3)
	adder1 : adder port map (N => COUNTER_OTPT, S => "0001", OTPT => ADDER1_OTPT);
	adder2 : adder port map (N => COUNTER_OTPT, S => "0010", OTPT => ADDER2_OTPT);
	adder3 : adder port map (N => COUNTER_OTPT, S => "0011", OTPT => ADDER3_OTPT);

	-- 4 instance of decodifier (3 bits to hex map)
	decodifier1 : decodifier port map (A => COUNTER_OTPT, OTPT => HEX3);
	decodifier2 : decodifier port map (A => ADDER1_OTPT, OTPT => HEX2);
	decodifier3 : decodifier port map (A => ADDER2_OTPT, OTPT => HEX1);
	decodifier4 : decodifier port map (A => ADDER3_OTPT, OTPT => HEX0);
	
	-- just for feedback (ledg show counter sequence, ledr(9) shows mux result)
	LEDG(0) <= COUNTER_OTPT(0);
	LEDG(1) <= COUNTER_OTPT(1);
	LEDG(2) <= COUNTER_OTPT(2);
	LEDG(3) <= COUNTER_OTPT(3);

	LEDR(9) <= MUX_OTPT;
end letter_arc;